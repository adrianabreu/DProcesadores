// first_nios2_system.v

// Generated using ACDS version 12.1sp1 243 at 2015.06.04.12:56:54

`timescale 1 ps / 1 ps
module first_nios2_system (
		inout  wire [15:0] sram_external_interface_DQ,         //     sram_external_interface.DQ
		output wire [17:0] sram_external_interface_ADDR,       //                            .ADDR
		output wire        sram_external_interface_LB_N,       //                            .LB_N
		output wire        sram_external_interface_UB_N,       //                            .UB_N
		output wire        sram_external_interface_CE_N,       //                            .CE_N
		output wire        sram_external_interface_OE_N,       //                            .OE_N
		output wire        sram_external_interface_WE_N,       //                            .WE_N
		output wire [7:0]  led_pio_external_connection_export, // led_pio_external_connection.export
		output wire [11:0] sdram_wire_addr,                    //                  sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                      //                            .ba
		output wire        sdram_wire_cas_n,                   //                            .cas_n
		output wire        sdram_wire_cke,                     //                            .cke
		output wire        sdram_wire_cs_n,                    //                            .cs_n
		inout  wire [15:0] sdram_wire_dq,                      //                            .dq
		output wire [1:0]  sdram_wire_dqm,                     //                            .dqm
		output wire        sdram_wire_ras_n,                   //                            .ras_n
		output wire        sdram_wire_we_n,                    //                            .we_n
		input  wire        reset_reset_n,                      //                       reset.reset_n
		input  wire        clk_clk,                            //                         clk.clk
		output wire        sdram_clk_clk                       //                   sdram_clk.clk
	);

	wire          clocks_sys_clk_clk;                                                                               // clocks:sys_clk -> [addr_router:clk, addr_router_001:clk, burst_adapter:clk, burst_adapter_001:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_003:clk, cpu:clk, cpu_data_master_translator:clk, cpu_data_master_translator_avalon_universal_master_0_agent:clk, cpu_instruction_master_translator:clk, cpu_instruction_master_translator_avalon_universal_master_0_agent:clk, cpu_jtag_debug_module_translator:clk, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, irq_mapper:clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, led_pio:clk, led_pio_s1_translator:clk, led_pio_s1_translator_avalon_universal_slave_0_agent:clk, led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, onchip_mem:clk, onchip_mem_s1_translator:clk, onchip_mem_s1_translator_avalon_universal_slave_0_agent:clk, onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, sdram:clk, sdram_s1_translator:clk, sdram_s1_translator_avalon_universal_slave_0_agent:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sram:clk, sram_avalon_sram_slave_translator:clk, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sys_clk_timer:clk, sys_clk_timer_s1_translator:clk, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:clk, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sysid:clock, sysid_control_slave_translator:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timestamp:clk, timestamp_s1_translator:clk, timestamp_s1_translator_avalon_universal_slave_0_agent:clk, timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk]
	wire          cpu_instruction_master_waitrequest;                                                               // cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	wire   [24:0] cpu_instruction_master_address;                                                                   // cpu:i_address -> cpu_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                      // cpu:i_read -> cpu_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                  // cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	wire          cpu_instruction_master_readdatavalid;                                                             // cpu_instruction_master_translator:av_readdatavalid -> cpu:i_readdatavalid
	wire          cpu_data_master_waitrequest;                                                                      // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                        // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire   [24:0] cpu_data_master_address;                                                                          // cpu:d_address -> cpu_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                            // cpu:d_write -> cpu_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                             // cpu:d_read -> cpu_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                         // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                                                      // cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	wire    [3:0] cpu_data_master_byteenable;                                                                       // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_jtag_debug_module_translator:av_chipselect -> cpu:jtag_debug_module_select
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_jtag_debug_module_translator:av_begintransfer -> cpu:jtag_debug_module_begintransfer
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	wire   [31:0] onchip_mem_s1_translator_avalon_anti_slave_0_writedata;                                           // onchip_mem_s1_translator:av_writedata -> onchip_mem:writedata
	wire   [12:0] onchip_mem_s1_translator_avalon_anti_slave_0_address;                                             // onchip_mem_s1_translator:av_address -> onchip_mem:address
	wire          onchip_mem_s1_translator_avalon_anti_slave_0_chipselect;                                          // onchip_mem_s1_translator:av_chipselect -> onchip_mem:chipselect
	wire          onchip_mem_s1_translator_avalon_anti_slave_0_clken;                                               // onchip_mem_s1_translator:av_clken -> onchip_mem:clken
	wire          onchip_mem_s1_translator_avalon_anti_slave_0_write;                                               // onchip_mem_s1_translator:av_write -> onchip_mem:write
	wire   [31:0] onchip_mem_s1_translator_avalon_anti_slave_0_readdata;                                            // onchip_mem:readdata -> onchip_mem_s1_translator:av_readdata
	wire    [3:0] onchip_mem_s1_translator_avalon_anti_slave_0_byteenable;                                          // onchip_mem_s1_translator:av_byteenable -> onchip_mem:byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                              // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [21:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                  // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                               // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                    // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                     // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                 // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                            // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                               // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                  // sram_avalon_sram_slave_translator:av_writedata -> sram:writedata
	wire   [17:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                    // sram_avalon_sram_slave_translator:av_address -> sram:address
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                      // sram_avalon_sram_slave_translator:av_write -> sram:write
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                       // sram_avalon_sram_slave_translator:av_read -> sram:read
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                   // sram:readdata -> sram_avalon_sram_slave_translator:av_readdata
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                              // sram:readdatavalid -> sram_avalon_sram_slave_translator:av_readdatavalid
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                 // sram_avalon_sram_slave_translator:av_byteenable -> sram:byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata;                                        // sys_clk_timer_s1_translator:av_writedata -> sys_clk_timer:writedata
	wire    [2:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_address;                                          // sys_clk_timer_s1_translator:av_address -> sys_clk_timer:address
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect;                                       // sys_clk_timer_s1_translator:av_chipselect -> sys_clk_timer:chipselect
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_write;                                            // sys_clk_timer_s1_translator:av_write -> sys_clk_timer:write_n
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata;                                         // sys_clk_timer:readdata -> sys_clk_timer_s1_translator:av_readdata
	wire    [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                       // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                      // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire   [31:0] led_pio_s1_translator_avalon_anti_slave_0_writedata;                                              // led_pio_s1_translator:av_writedata -> led_pio:writedata
	wire    [1:0] led_pio_s1_translator_avalon_anti_slave_0_address;                                                // led_pio_s1_translator:av_address -> led_pio:address
	wire          led_pio_s1_translator_avalon_anti_slave_0_chipselect;                                             // led_pio_s1_translator:av_chipselect -> led_pio:chipselect
	wire          led_pio_s1_translator_avalon_anti_slave_0_write;                                                  // led_pio_s1_translator:av_write -> led_pio:write_n
	wire   [31:0] led_pio_s1_translator_avalon_anti_slave_0_readdata;                                               // led_pio:readdata -> led_pio_s1_translator:av_readdata
	wire   [15:0] timestamp_s1_translator_avalon_anti_slave_0_writedata;                                            // timestamp_s1_translator:av_writedata -> timestamp:writedata
	wire    [3:0] timestamp_s1_translator_avalon_anti_slave_0_address;                                              // timestamp_s1_translator:av_address -> timestamp:address
	wire          timestamp_s1_translator_avalon_anti_slave_0_chipselect;                                           // timestamp_s1_translator:av_chipselect -> timestamp:chipselect
	wire          timestamp_s1_translator_avalon_anti_slave_0_write;                                                // timestamp_s1_translator:av_write -> timestamp:write_n
	wire   [15:0] timestamp_s1_translator_avalon_anti_slave_0_readdata;                                             // timestamp:readdata -> timestamp_s1_translator:av_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [24:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [24:0] cpu_data_master_translator_avalon_universal_master_0_address;                                     // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                       // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                        // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	wire   [24:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // onchip_mem_s1_translator:uav_waitrequest -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_mem_s1_translator:uav_burstcount
	wire   [31:0] onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_mem_s1_translator:uav_writedata
	wire   [24:0] onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_mem_s1_translator:uav_address
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_mem_s1_translator:uav_write
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_mem_s1_translator:uav_lock
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_mem_s1_translator:uav_read
	wire   [31:0] onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // onchip_mem_s1_translator:uav_readdata -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // onchip_mem_s1_translator:uav_readdatavalid -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_mem_s1_translator:uav_debugaccess
	wire    [3:0] onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_mem_s1_translator:uav_byteenable
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [24:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // sram_avalon_sram_slave_translator:uav_waitrequest -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_avalon_sram_slave_translator:uav_burstcount
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                    // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_avalon_sram_slave_translator:uav_writedata
	wire   [24:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                      // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> sram_avalon_sram_slave_translator:uav_address
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                        // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> sram_avalon_sram_slave_translator:uav_write
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                         // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sram_avalon_sram_slave_translator:uav_lock
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                         // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> sram_avalon_sram_slave_translator:uav_read
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                     // sram_avalon_sram_slave_translator:uav_readdata -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // sram_avalon_sram_slave_translator:uav_readdatavalid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_avalon_sram_slave_translator:uav_debugaccess
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_avalon_sram_slave_translator:uav_byteenable
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                  // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire   [24:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // sys_clk_timer_s1_translator:uav_waitrequest -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sys_clk_timer_s1_translator:uav_burstcount
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sys_clk_timer_s1_translator:uav_writedata
	wire   [24:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> sys_clk_timer_s1_translator:uav_address
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> sys_clk_timer_s1_translator:uav_write
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sys_clk_timer_s1_translator:uav_lock
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> sys_clk_timer_s1_translator:uav_read
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // sys_clk_timer_s1_translator:uav_readdata -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // sys_clk_timer_s1_translator:uav_readdatavalid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sys_clk_timer_s1_translator:uav_debugaccess
	wire    [3:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sys_clk_timer_s1_translator:uav_byteenable
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire   [24:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // led_pio_s1_translator:uav_waitrequest -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_pio_s1_translator:uav_burstcount
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_pio_s1_translator:uav_writedata
	wire   [24:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_pio_s1_translator:uav_address
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_pio_s1_translator:uav_write
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_pio_s1_translator:uav_lock
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_pio_s1_translator:uav_read
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // led_pio_s1_translator:uav_readdata -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // led_pio_s1_translator:uav_readdatavalid -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_pio_s1_translator:uav_debugaccess
	wire    [3:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_pio_s1_translator:uav_byteenable
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // timestamp_s1_translator:uav_waitrequest -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timestamp_s1_translator:uav_burstcount
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timestamp_s1_translator:uav_writedata
	wire   [24:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_address -> timestamp_s1_translator:uav_address
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_write -> timestamp_s1_translator:uav_write
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timestamp_s1_translator:uav_lock
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_read -> timestamp_s1_translator:uav_read
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // timestamp_s1_translator:uav_readdata -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // timestamp_s1_translator:uav_readdatavalid -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timestamp_s1_translator:uav_debugaccess
	wire    [3:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timestamp_s1_translator:uav_byteenable
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire   [99:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire   [99:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_001:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire   [99:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [99:0] onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // onchip_mem_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_001:sink_ready -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [81:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_002:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                        // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire   [81:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                         // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_003:sink_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire   [99:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_004:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire   [99:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_005:sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire   [99:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_006:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [99:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_007:sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire   [99:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_008:sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                      // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                            // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                    // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire   [99:0] addr_router_src_data;                                                                             // addr_router:src_data -> limiter:cmd_sink_data
	wire    [8:0] addr_router_src_channel;                                                                          // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                            // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                      // limiter:rsp_src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                            // limiter:rsp_src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                    // limiter:rsp_src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [99:0] limiter_rsp_src_data;                                                                             // limiter:rsp_src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [8:0] limiter_rsp_src_channel;                                                                          // limiter:rsp_src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                            // cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                // burst_adapter:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                      // burst_adapter:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                              // burst_adapter:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] burst_adapter_source0_data;                                                                       // burst_adapter:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                      // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [8:0] burst_adapter_source0_channel;                                                                    // burst_adapter:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                            // burst_adapter_001:source0_endofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                  // burst_adapter_001:source0_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                          // burst_adapter_001:source0_startofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] burst_adapter_001_source0_data;                                                                   // burst_adapter_001:source0_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                  // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire    [8:0] burst_adapter_001_source0_channel;                                                                // burst_adapter_001:source0_channel -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                   // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, irq_mapper:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_pio:reset_n, led_pio_s1_translator:reset, led_pio_s1_translator_avalon_universal_slave_0_agent:reset, led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, onchip_mem:reset, onchip_mem_s1_translator:reset, onchip_mem_s1_translator_avalon_universal_slave_0_agent:reset, onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sram:reset, sram_avalon_sram_slave_translator:reset, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sys_clk_timer:reset_n, sys_clk_timer_s1_translator:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timestamp:reset_n, timestamp_s1_translator:reset, timestamp_s1_translator_avalon_universal_slave_0_agent:reset, timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire          rst_controller_001_reset_out_reset;                                                               // rst_controller_001:reset_out -> clocks:reset
	wire          cmd_xbar_demux_src0_endofpacket;                                                                  // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                        // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire   [99:0] cmd_xbar_demux_src0_data;                                                                         // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire    [8:0] cmd_xbar_demux_src0_channel;                                                                      // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                        // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                  // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                        // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire   [99:0] cmd_xbar_demux_src1_data;                                                                         // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire    [8:0] cmd_xbar_demux_src1_channel;                                                                      // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                        // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                  // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                        // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire   [99:0] cmd_xbar_demux_src2_data;                                                                         // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire    [8:0] cmd_xbar_demux_src2_channel;                                                                      // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                        // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                  // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                        // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire   [99:0] cmd_xbar_demux_src3_data;                                                                         // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire    [8:0] cmd_xbar_demux_src3_channel;                                                                      // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                        // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                              // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                    // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                            // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src0_data;                                                                     // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire    [8:0] cmd_xbar_demux_001_src0_channel;                                                                  // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                    // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                              // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                    // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                            // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src1_data;                                                                     // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire    [8:0] cmd_xbar_demux_001_src1_channel;                                                                  // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                    // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                              // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                    // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                            // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src2_data;                                                                     // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire    [8:0] cmd_xbar_demux_001_src2_channel;                                                                  // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                    // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                              // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                    // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                            // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src3_data;                                                                     // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire    [8:0] cmd_xbar_demux_001_src3_channel;                                                                  // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                    // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                              // cmd_xbar_demux_001:src4_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                    // cmd_xbar_demux_001:src4_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                            // cmd_xbar_demux_001:src4_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src4_data;                                                                     // cmd_xbar_demux_001:src4_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_demux_001_src4_channel;                                                                  // cmd_xbar_demux_001:src4_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                              // cmd_xbar_demux_001:src5_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                    // cmd_xbar_demux_001:src5_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                            // cmd_xbar_demux_001:src5_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src5_data;                                                                     // cmd_xbar_demux_001:src5_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_demux_001_src5_channel;                                                                  // cmd_xbar_demux_001:src5_channel -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                              // cmd_xbar_demux_001:src6_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                    // cmd_xbar_demux_001:src6_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                            // cmd_xbar_demux_001:src6_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src6_data;                                                                     // cmd_xbar_demux_001:src6_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_demux_001_src6_channel;                                                                  // cmd_xbar_demux_001:src6_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                              // cmd_xbar_demux_001:src7_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                    // cmd_xbar_demux_001:src7_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                            // cmd_xbar_demux_001:src7_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src7_data;                                                                     // cmd_xbar_demux_001:src7_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_demux_001_src7_channel;                                                                  // cmd_xbar_demux_001:src7_channel -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                              // cmd_xbar_demux_001:src8_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                    // cmd_xbar_demux_001:src8_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                            // cmd_xbar_demux_001:src8_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src8_data;                                                                     // cmd_xbar_demux_001:src8_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_demux_001_src8_channel;                                                                  // cmd_xbar_demux_001:src8_channel -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                  // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                        // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire   [99:0] rsp_xbar_demux_src0_data;                                                                         // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [8:0] rsp_xbar_demux_src0_channel;                                                                      // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                        // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                  // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                        // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire   [99:0] rsp_xbar_demux_src1_data;                                                                         // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire    [8:0] rsp_xbar_demux_src1_channel;                                                                      // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                        // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                              // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                    // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                            // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire   [99:0] rsp_xbar_demux_001_src0_data;                                                                     // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [8:0] rsp_xbar_demux_001_src0_channel;                                                                  // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                    // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                              // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                    // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                            // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire   [99:0] rsp_xbar_demux_001_src1_data;                                                                     // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire    [8:0] rsp_xbar_demux_001_src1_channel;                                                                  // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                    // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                              // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                    // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                            // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire   [99:0] rsp_xbar_demux_002_src0_data;                                                                     // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [8:0] rsp_xbar_demux_002_src0_channel;                                                                  // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                    // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                              // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                    // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                            // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire   [99:0] rsp_xbar_demux_002_src1_data;                                                                     // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire    [8:0] rsp_xbar_demux_002_src1_channel;                                                                  // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                    // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                              // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                    // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                            // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire   [99:0] rsp_xbar_demux_003_src0_data;                                                                     // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire    [8:0] rsp_xbar_demux_003_src0_channel;                                                                  // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                    // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                              // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                    // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                            // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire   [99:0] rsp_xbar_demux_003_src1_data;                                                                     // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire    [8:0] rsp_xbar_demux_003_src1_channel;                                                                  // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                    // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                              // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                    // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                            // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire   [99:0] rsp_xbar_demux_004_src0_data;                                                                     // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire    [8:0] rsp_xbar_demux_004_src0_channel;                                                                  // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                    // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                              // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                    // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                            // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire   [99:0] rsp_xbar_demux_005_src0_data;                                                                     // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire    [8:0] rsp_xbar_demux_005_src0_channel;                                                                  // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                    // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                              // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                    // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                            // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire   [99:0] rsp_xbar_demux_006_src0_data;                                                                     // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire    [8:0] rsp_xbar_demux_006_src0_channel;                                                                  // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                    // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                              // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                    // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                            // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire   [99:0] rsp_xbar_demux_007_src0_data;                                                                     // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire    [8:0] rsp_xbar_demux_007_src0_channel;                                                                  // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                    // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                              // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                    // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                            // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire   [99:0] rsp_xbar_demux_008_src0_data;                                                                     // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire    [8:0] rsp_xbar_demux_008_src0_channel;                                                                  // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                    // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                      // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                    // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire   [99:0] limiter_cmd_src_data;                                                                             // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire    [8:0] limiter_cmd_src_channel;                                                                          // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                            // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                     // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                           // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                   // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire   [99:0] rsp_xbar_mux_src_data;                                                                            // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire    [8:0] rsp_xbar_mux_src_channel;                                                                         // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                           // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                  // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                        // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire   [99:0] addr_router_001_src_data;                                                                         // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [8:0] addr_router_001_src_channel;                                                                      // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                        // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                 // rsp_xbar_mux_001:src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                       // rsp_xbar_mux_001:src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                               // rsp_xbar_mux_001:src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [99:0] rsp_xbar_mux_001_src_data;                                                                        // rsp_xbar_mux_001:src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [8:0] rsp_xbar_mux_001_src_channel;                                                                     // rsp_xbar_mux_001:src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                       // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                     // cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                           // cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                   // cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_mux_src_data;                                                                            // cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_mux_src_channel;                                                                         // cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                        // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                              // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                      // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire   [99:0] id_router_src_data;                                                                               // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [8:0] id_router_src_channel;                                                                            // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                              // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                 // cmd_xbar_mux_001:src_endofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                       // cmd_xbar_mux_001:src_valid -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                               // cmd_xbar_mux_001:src_startofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_mux_001_src_data;                                                                        // cmd_xbar_mux_001:src_data -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_mux_001_src_channel;                                                                     // cmd_xbar_mux_001:src_channel -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                       // onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                    // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                          // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                  // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire   [99:0] id_router_001_src_data;                                                                           // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [8:0] id_router_001_src_channel;                                                                        // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                          // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                    // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                          // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                  // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire   [99:0] id_router_004_src_data;                                                                           // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [8:0] id_router_004_src_channel;                                                                        // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                          // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                    // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                          // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                  // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire   [99:0] id_router_005_src_data;                                                                           // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire    [8:0] id_router_005_src_channel;                                                                        // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                          // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                    // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                          // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                  // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire   [99:0] id_router_006_src_data;                                                                           // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire    [8:0] id_router_006_src_channel;                                                                        // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                          // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                    // led_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                    // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                          // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                  // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [99:0] id_router_007_src_data;                                                                           // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire    [8:0] id_router_007_src_channel;                                                                        // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                          // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                    // timestamp_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                    // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                          // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                  // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [99:0] id_router_008_src_data;                                                                           // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire    [8:0] id_router_008_src_channel;                                                                        // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                          // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                 // cmd_xbar_mux_002:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                       // cmd_xbar_mux_002:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                               // cmd_xbar_mux_002:src_startofpacket -> width_adapter:in_startofpacket
	wire   [99:0] cmd_xbar_mux_002_src_data;                                                                        // cmd_xbar_mux_002:src_data -> width_adapter:in_data
	wire    [8:0] cmd_xbar_mux_002_src_channel;                                                                     // cmd_xbar_mux_002:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                       // width_adapter:in_ready -> cmd_xbar_mux_002:src_ready
	wire          width_adapter_src_endofpacket;                                                                    // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                          // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                  // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [81:0] width_adapter_src_data;                                                                           // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                          // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire    [8:0] width_adapter_src_channel;                                                                        // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_002_src_endofpacket;                                                                    // id_router_002:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_002_src_valid;                                                                          // id_router_002:src_valid -> width_adapter_001:in_valid
	wire          id_router_002_src_startofpacket;                                                                  // id_router_002:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [81:0] id_router_002_src_data;                                                                           // id_router_002:src_data -> width_adapter_001:in_data
	wire    [8:0] id_router_002_src_channel;                                                                        // id_router_002:src_channel -> width_adapter_001:in_channel
	wire          id_router_002_src_ready;                                                                          // width_adapter_001:in_ready -> id_router_002:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                // width_adapter_001:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                      // width_adapter_001:out_valid -> rsp_xbar_demux_002:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                              // width_adapter_001:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire   [99:0] width_adapter_001_src_data;                                                                       // width_adapter_001:out_data -> rsp_xbar_demux_002:sink_data
	wire          width_adapter_001_src_ready;                                                                      // rsp_xbar_demux_002:sink_ready -> width_adapter_001:out_ready
	wire    [8:0] width_adapter_001_src_channel;                                                                    // width_adapter_001:out_channel -> rsp_xbar_demux_002:sink_channel
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                 // cmd_xbar_mux_003:src_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                       // cmd_xbar_mux_003:src_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                               // cmd_xbar_mux_003:src_startofpacket -> width_adapter_002:in_startofpacket
	wire   [99:0] cmd_xbar_mux_003_src_data;                                                                        // cmd_xbar_mux_003:src_data -> width_adapter_002:in_data
	wire    [8:0] cmd_xbar_mux_003_src_channel;                                                                     // cmd_xbar_mux_003:src_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                       // width_adapter_002:in_ready -> cmd_xbar_mux_003:src_ready
	wire          width_adapter_002_src_endofpacket;                                                                // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                      // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                              // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [81:0] width_adapter_002_src_data;                                                                       // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire          width_adapter_002_src_ready;                                                                      // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire    [8:0] width_adapter_002_src_channel;                                                                    // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          id_router_003_src_endofpacket;                                                                    // id_router_003:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_003_src_valid;                                                                          // id_router_003:src_valid -> width_adapter_003:in_valid
	wire          id_router_003_src_startofpacket;                                                                  // id_router_003:src_startofpacket -> width_adapter_003:in_startofpacket
	wire   [81:0] id_router_003_src_data;                                                                           // id_router_003:src_data -> width_adapter_003:in_data
	wire    [8:0] id_router_003_src_channel;                                                                        // id_router_003:src_channel -> width_adapter_003:in_channel
	wire          id_router_003_src_ready;                                                                          // width_adapter_003:in_ready -> id_router_003:src_ready
	wire          width_adapter_003_src_endofpacket;                                                                // width_adapter_003:out_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                                      // width_adapter_003:out_valid -> rsp_xbar_demux_003:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                              // width_adapter_003:out_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire   [99:0] width_adapter_003_src_data;                                                                       // width_adapter_003:out_data -> rsp_xbar_demux_003:sink_data
	wire          width_adapter_003_src_ready;                                                                      // rsp_xbar_demux_003:sink_ready -> width_adapter_003:out_ready
	wire    [8:0] width_adapter_003_src_channel;                                                                    // width_adapter_003:out_channel -> rsp_xbar_demux_003:sink_channel
	wire    [8:0] limiter_cmd_valid_data;                                                                           // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                         // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                         // sys_clk_timer:irq -> irq_mapper:receiver1_irq
	wire   [31:0] cpu_d_irq_irq;                                                                                    // irq_mapper:sender_irq -> cpu:d_irq

	first_nios2_system_onchip_mem onchip_mem (
		.clk        (clocks_sys_clk_clk),                                      //   clk1.clk
		.address    (onchip_mem_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_mem_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_mem_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_mem_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_mem_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_mem_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_mem_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                           // reset1.reset
	);

	first_nios2_system_cpu cpu (
		.clk                                   (clocks_sys_clk_clk),                                                 //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                    //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	first_nios2_system_jtag_uart jtag_uart (
		.clk            (clocks_sys_clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	first_nios2_system_sys_clk_timer sys_clk_timer (
		.clk        (clocks_sys_clk_clk),                                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                            // reset.reset_n
		.address    (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~sys_clk_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                                    //   irq.irq
	);

	first_nios2_system_sysid sysid (
		.clock    (clocks_sys_clk_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                             //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	first_nios2_system_led_pio led_pio (
		.clk        (clocks_sys_clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (led_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_pio_external_connection_export)                    // external_connection.export
	);

	first_nios2_system_sdram sdram (
		.clk            (clocks_sys_clk_clk),                                    //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                       // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	first_nios2_system_clocks clocks (
		.CLOCK_50    (clk_clk),                            //       clk_in_primary.clk
		.reset       (rst_controller_001_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (clocks_sys_clk_clk),                 //              sys_clk.clk
		.sys_reset_n (),                                   //        sys_clk_reset.reset_n
		.SDRAM_CLK   (sdram_clk_clk)                       //            sdram_clk.clk
	);

	first_nios2_system_sram sram (
		.clk           (clocks_sys_clk_clk),                                                  //        clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                      //  clock_reset_reset.reset
		.SRAM_DQ       (sram_external_interface_DQ),                                          // external_interface.export
		.SRAM_ADDR     (sram_external_interface_ADDR),                                        //                   .export
		.SRAM_LB_N     (sram_external_interface_LB_N),                                        //                   .export
		.SRAM_UB_N     (sram_external_interface_UB_N),                                        //                   .export
		.SRAM_CE_N     (sram_external_interface_CE_N),                                        //                   .export
		.SRAM_OE_N     (sram_external_interface_OE_N),                                        //                   .export
		.SRAM_WE_N     (sram_external_interface_WE_N),                                        //                   .export
		.address       (sram_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (sram_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (sram_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	first_nios2_system_timestamp timestamp (
		.clk        (clocks_sys_clk_clk),                                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        // reset.reset_n
		.address    (timestamp_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timestamp_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timestamp_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timestamp_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timestamp_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        ()                                                        //   irq.irq
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                   (clocks_sys_clk_clk),                                                        //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address           (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                      //               (terminated)
		.av_byteenable         (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_write              (1'b0),                                                                      //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.av_debugaccess        (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                   (clocks_sys_clk_clk),                                                 //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address           (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_data_master_read),                                               //                          .read
		.av_readdata           (cpu_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_data_master_write),                                              //                          .write
		.av_writedata          (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_readdatavalid      (),                                                                   //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                   (clocks_sys_clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_mem_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_mem_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_mem_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_mem_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_mem_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_mem_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_mem_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_mem_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sram_avalon_sram_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sram_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sram_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sram_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_chipselect         (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sys_clk_timer_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sys_clk_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_writedata          (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_pio_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                    //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (led_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (led_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (led_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (led_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (led_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timestamp_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timestamp_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timestamp_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timestamp_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timestamp_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timestamp_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_BEGIN_BURST           (80),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.PKT_BURST_TYPE_H          (77),
		.PKT_BURST_TYPE_L          (76),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (86),
		.PKT_THREAD_ID_H           (90),
		.PKT_THREAD_ID_L           (90),
		.PKT_CACHE_H               (97),
		.PKT_CACHE_L               (94),
		.PKT_DATA_SIDEBAND_H       (79),
		.PKT_DATA_SIDEBAND_L       (79),
		.PKT_QOS_H                 (81),
		.PKT_QOS_L                 (81),
		.PKT_ADDR_SIDEBAND_H       (78),
		.PKT_ADDR_SIDEBAND_L       (78),
		.ST_DATA_W                 (100),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clocks_sys_clk_clk),                                                                 //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address       (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                              //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                               //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                               //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_BEGIN_BURST           (80),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.PKT_BURST_TYPE_H          (77),
		.PKT_BURST_TYPE_L          (76),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (86),
		.PKT_THREAD_ID_H           (90),
		.PKT_THREAD_ID_L           (90),
		.PKT_CACHE_H               (97),
		.PKT_CACHE_L               (94),
		.PKT_DATA_SIDEBAND_H       (79),
		.PKT_DATA_SIDEBAND_L       (79),
		.PKT_QOS_H                 (81),
		.PKT_QOS_L                 (81),
		.PKT_ADDR_SIDEBAND_H       (78),
		.PKT_ADDR_SIDEBAND_L       (78),
		.ST_DATA_W                 (100),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clocks_sys_clk_clk),                                                          //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address       (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                  //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                   //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                          //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                            //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                   //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_mem_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                       //                .channel
		.rf_sink_ready           (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (62),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                   //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                   //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                    //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                             //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                 //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (62),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                             //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                             //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                              //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                       //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                           //                .channel
		.rf_sink_ready           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                       //                .channel
		.rf_sink_ready           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) led_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                 //                .channel
		.rf_sink_ready           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timestamp_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                   //                .channel
		.rf_sink_ready           (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	first_nios2_system_addr_router addr_router (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	first_nios2_system_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                              //          .endofpacket
	);

	first_nios2_system_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	first_nios2_system_id_router id_router_001 (
		.sink_ready         (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                  //       src.ready
		.src_valid          (id_router_001_src_valid),                                                  //          .valid
		.src_data           (id_router_001_src_data),                                                   //          .data
		.src_channel        (id_router_001_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                             //          .endofpacket
	);

	first_nios2_system_id_router_002 id_router_002 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                             //       src.ready
		.src_valid          (id_router_002_src_valid),                                             //          .valid
		.src_data           (id_router_002_src_data),                                              //          .data
		.src_channel        (id_router_002_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                        //          .endofpacket
	);

	first_nios2_system_id_router_002 id_router_003 (
		.sink_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                           //       src.ready
		.src_valid          (id_router_003_src_valid),                                                           //          .valid
		.src_data           (id_router_003_src_data),                                                            //          .data
		.src_channel        (id_router_003_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                      //          .endofpacket
	);

	first_nios2_system_id_router_004 id_router_004 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                //          .valid
		.src_data           (id_router_004_src_data),                                                                 //          .data
		.src_channel        (id_router_004_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                           //          .endofpacket
	);

	first_nios2_system_id_router_004 id_router_005 (
		.sink_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                     //       src.ready
		.src_valid          (id_router_005_src_valid),                                                     //          .valid
		.src_data           (id_router_005_src_data),                                                      //          .data
		.src_channel        (id_router_005_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                //          .endofpacket
	);

	first_nios2_system_id_router_004 id_router_006 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                        //       src.ready
		.src_valid          (id_router_006_src_valid),                                                        //          .valid
		.src_data           (id_router_006_src_data),                                                         //          .data
		.src_channel        (id_router_006_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                   //          .endofpacket
	);

	first_nios2_system_id_router_004 id_router_007 (
		.sink_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                               //       src.ready
		.src_valid          (id_router_007_src_valid),                                               //          .valid
		.src_data           (id_router_007_src_data),                                                //          .data
		.src_channel        (id_router_007_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                          //          .endofpacket
	);

	first_nios2_system_id_router_004 id_router_008 (
		.sink_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                 //       src.ready
		.src_valid          (id_router_008_src_valid),                                                 //          .valid
		.src_data           (id_router_008_src_data),                                                  //          .data
		.src_channel        (id_router_008_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                            //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (86),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (100),
		.ST_CHANNEL_W              (9),
		.VALID_WIDTH               (9),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clocks_sys_clk_clk),             //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (62),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.PKT_BURST_TYPE_H          (59),
		.PKT_BURST_TYPE_L          (58),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (9),
		.OUT_BYTE_CNT_H            (50),
		.OUT_BURSTWRAP_H           (54),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clocks_sys_clk_clk),                  //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (62),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.PKT_BURST_TYPE_H          (59),
		.PKT_BURST_TYPE_L          (58),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (9),
		.OUT_BYTE_CNT_H            (50),
		.OUT_BURSTWRAP_H           (54),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clocks_sys_clk_clk),             //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	first_nios2_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clocks_sys_clk_clk),                //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)    //           .endofpacket
	);

	first_nios2_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //          .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),         //      src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),         //          .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),          //          .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),       //          .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //          .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),         //      src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket),   //          .endofpacket
		.src8_ready         (cmd_xbar_demux_001_src8_ready),         //      src8.ready
		.src8_valid         (cmd_xbar_demux_001_src8_valid),         //          .valid
		.src8_data          (cmd_xbar_demux_001_src8_data),          //          .data
		.src8_channel       (cmd_xbar_demux_001_src8_channel),       //          .channel
		.src8_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_001_src8_endofpacket)    //          .endofpacket
	);

	first_nios2_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	first_nios2_system_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	first_nios2_system_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	first_nios2_system_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	first_nios2_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clocks_sys_clk_clk),                //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	first_nios2_system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	first_nios2_system_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	first_nios2_system_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	first_nios2_system_rsp_xbar_demux_004 rsp_xbar_demux_004 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	first_nios2_system_rsp_xbar_demux_004 rsp_xbar_demux_005 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	first_nios2_system_rsp_xbar_demux_004 rsp_xbar_demux_006 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	first_nios2_system_rsp_xbar_demux_004 rsp_xbar_demux_007 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	first_nios2_system_rsp_xbar_demux_004 rsp_xbar_demux_008 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	first_nios2_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	first_nios2_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready         (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (69),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (72),
		.IN_PKT_BURSTWRAP_L            (70),
		.IN_PKT_BURST_SIZE_H           (75),
		.IN_PKT_BURST_SIZE_L           (73),
		.IN_PKT_RESPONSE_STATUS_H      (99),
		.IN_PKT_RESPONSE_STATUS_L      (98),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (77),
		.IN_PKT_BURST_TYPE_L           (76),
		.IN_ST_DATA_W                  (100),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (51),
		.OUT_PKT_BYTE_CNT_L            (49),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_PKT_BURST_SIZE_H          (57),
		.OUT_PKT_BURST_SIZE_L          (55),
		.OUT_PKT_RESPONSE_STATUS_H     (81),
		.OUT_PKT_RESPONSE_STATUS_L     (80),
		.OUT_PKT_TRANS_EXCLUSIVE       (48),
		.OUT_PKT_BURST_TYPE_H          (59),
		.OUT_PKT_BURST_TYPE_L          (58),
		.OUT_ST_DATA_W                 (82),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (clocks_sys_clk_clk),                 //       clk.clk
		.reset                (rst_controller_reset_out_reset),     // clk_reset.reset
		.in_valid             (cmd_xbar_mux_002_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_002_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_002_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_002_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_002_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (51),
		.IN_PKT_BYTE_CNT_L             (49),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (54),
		.IN_PKT_BURSTWRAP_L            (52),
		.IN_PKT_BURST_SIZE_H           (57),
		.IN_PKT_BURST_SIZE_L           (55),
		.IN_PKT_RESPONSE_STATUS_H      (81),
		.IN_PKT_RESPONSE_STATUS_L      (80),
		.IN_PKT_TRANS_EXCLUSIVE        (48),
		.IN_PKT_BURST_TYPE_H           (59),
		.IN_PKT_BURST_TYPE_L           (58),
		.IN_ST_DATA_W                  (82),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (69),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (75),
		.OUT_PKT_BURST_SIZE_L          (73),
		.OUT_PKT_RESPONSE_STATUS_H     (99),
		.OUT_PKT_RESPONSE_STATUS_L     (98),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (77),
		.OUT_PKT_BURST_TYPE_L          (76),
		.OUT_ST_DATA_W                 (100),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (clocks_sys_clk_clk),                  //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_002_src_valid),             //      sink.valid
		.in_channel           (id_router_002_src_channel),           //          .channel
		.in_startofpacket     (id_router_002_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_002_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_002_src_ready),             //          .ready
		.in_data              (id_router_002_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (69),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (72),
		.IN_PKT_BURSTWRAP_L            (70),
		.IN_PKT_BURST_SIZE_H           (75),
		.IN_PKT_BURST_SIZE_L           (73),
		.IN_PKT_RESPONSE_STATUS_H      (99),
		.IN_PKT_RESPONSE_STATUS_L      (98),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (77),
		.IN_PKT_BURST_TYPE_L           (76),
		.IN_ST_DATA_W                  (100),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (51),
		.OUT_PKT_BYTE_CNT_L            (49),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_PKT_BURST_SIZE_H          (57),
		.OUT_PKT_BURST_SIZE_L          (55),
		.OUT_PKT_RESPONSE_STATUS_H     (81),
		.OUT_PKT_RESPONSE_STATUS_L     (80),
		.OUT_PKT_TRANS_EXCLUSIVE       (48),
		.OUT_PKT_BURST_TYPE_H          (59),
		.OUT_PKT_BURST_TYPE_L          (58),
		.OUT_ST_DATA_W                 (82),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk                  (clocks_sys_clk_clk),                  //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_mux_003_src_valid),          //      sink.valid
		.in_channel           (cmd_xbar_mux_003_src_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_mux_003_src_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_003_src_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_mux_003_src_ready),          //          .ready
		.in_data              (cmd_xbar_mux_003_src_data),           //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_002_src_data),          //          .data
		.out_channel          (width_adapter_002_src_channel),       //          .channel
		.out_valid            (width_adapter_002_src_valid),         //          .valid
		.out_ready            (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (51),
		.IN_PKT_BYTE_CNT_L             (49),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (54),
		.IN_PKT_BURSTWRAP_L            (52),
		.IN_PKT_BURST_SIZE_H           (57),
		.IN_PKT_BURST_SIZE_L           (55),
		.IN_PKT_RESPONSE_STATUS_H      (81),
		.IN_PKT_RESPONSE_STATUS_L      (80),
		.IN_PKT_TRANS_EXCLUSIVE        (48),
		.IN_PKT_BURST_TYPE_H           (59),
		.IN_PKT_BURST_TYPE_L           (58),
		.IN_ST_DATA_W                  (82),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (69),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (75),
		.OUT_PKT_BURST_SIZE_L          (73),
		.OUT_PKT_RESPONSE_STATUS_H     (99),
		.OUT_PKT_RESPONSE_STATUS_L     (98),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (77),
		.OUT_PKT_BURST_TYPE_L          (76),
		.OUT_ST_DATA_W                 (100),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_003 (
		.clk                  (clocks_sys_clk_clk),                  //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_003_src_valid),             //      sink.valid
		.in_channel           (id_router_003_src_channel),           //          .channel
		.in_startofpacket     (id_router_003_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_003_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_003_src_ready),             //          .ready
		.in_data              (id_router_003_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	first_nios2_system_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

endmodule
