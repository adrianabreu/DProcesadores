module ModuloSonido(input clk,
							output reg enable,
							input reset, short, long,
							output wire[51:0] sonido
							);
	reg[51:0] frecuencia;
	assign sonido= frecuencia;
	reg still;

	always@(clk)
		begin0
			if (short)
				begin
					enable <= 1;
					frecuencia <=  32000;
				end
			else
				begin
				if (long)
					begin
						enable <= 1;
						still <= 1;
						frecuencia <=  32000;
					end
				else
					begin
					if(still)
						begin
							still <= 0;
							enable <= 1;
							frecuencia <=  32000;
						end
					else
						begin
							enable <= 0;
							frecuencia <=  0;
						end
					end
				end
		end
endmodule
